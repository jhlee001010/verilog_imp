module vending_machine_controller(
    input clk;
    input reset;
    
    input Ba;
    input Bb;
    input Bc;
    
    input Sc;
    input Sp;



);

