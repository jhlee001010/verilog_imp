module tl_controller (


);